** Profile: "SCHEMATIC1-Practica 1-1"  [ C:\Users\uriel\Desktop\Practica 1\Practica 1.1\practica 1-1-pspicefiles\schematic1\practica 1-1.sim ] 

** Creating circuit file "Practica 1-1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN 50u 40m 0 50u 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
